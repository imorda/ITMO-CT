`include "cpu_test.v"